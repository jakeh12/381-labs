-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
-------------------------------------------------------------------------------
entity mips is
  
  port (
    i_clk : in std_logic;
    i_rst : in std_logic);

end entity mips;
-------------------------------------------------------------------------------
architecture mixed of mips is

begin  -- architecture mixed

  

  -----------------------------------------------------------------------------
  -- Main Control
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  -- PC and Instruction Fetch
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  -- Instruction Memory
  -----------------------------------------------------------------------------


  
  -----------------------------------------------------------------------------
  -- Register File
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  -- ALU Control
  -----------------------------------------------------------------------------


  -----------------------------------------------------------------------------
  -- ALU
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  -- Branch Control
  -----------------------------------------------------------------------------


  -----------------------------------------------------------------------------
  -- Data Memory
  -----------------------------------------------------------------------------

  
end architecture mixed;
-------------------------------------------------------------------------------
