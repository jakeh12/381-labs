-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
-------------------------------------------------------------------------------
entity mips_multiplier is
  
  port (
    i_A : in  std_logic_vector (31 downto 0);   -- multiplicant
    i_B : in  std_logic_vector (31 downto 0);   -- multiplier
    i_O : out std_logic_vector (31 downto 0));  -- product

end entity mips_multiplier;
-------------------------------------------------------------------------------
architecture mixed of mips_multiplier is

  
  
begin  -- architecture mixed

  

end architecture mixed;
-------------------------------------------------------------------------------
