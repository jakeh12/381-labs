library ieee;
use ieee.std_logic_1164.all;

entity decoder5to32 is
  port(i_X : in std_logic_vector(4 downto 0);     -- raw value
       i_En : in std_logic;
       o_Y : out std_logic_vector(31 downto 0));   -- decoded value
end decoder5to32;

architecture dataflow of decoder5to32 is

	signal s_Y : std_logic_vector(31 downto 0) := (others => '0');

begin

	o_Y <= s_Y when i_En = '1' else (others => '0');

	with i_X select
		s_Y <= "00000000000000000000000000000001" when "00000", -- 00
		       "00000000000000000000000000000010" when "00001", -- 01
		       "00000000000000000000000000000100" when "00010", -- 02
		       "00000000000000000000000000001000" when "00011", -- 03
		       "00000000000000000000000000010000" when "00100", -- 04
		       "00000000000000000000000000100000" when "00101", -- 05
		       "00000000000000000000000001000000" when "00110", -- 06
		       "00000000000000000000000010000000" when "00111", -- 07
		       "00000000000000000000000100000000" when "01000", -- 08
		       "00000000000000000000001000000000" when "01001", -- 09
		       "00000000000000000000010000000000" when "01010", -- 0A
		       "00000000000000000000100000000000" when "01011", -- 0B
		       "00000000000000000001000000000000" when "01100", -- 0C
		       "00000000000000000010000000000000" when "01101", -- 0D
		       "00000000000000000100000000000000" when "01110", -- 0E
		       "00000000000000001000000000000000" when "01111", -- 0F
		       "00000000000000010000000000000000" when "10000", -- 10
		       "00000000000000100000000000000000" when "10001", -- 11
		       "00000000000001000000000000000000" when "10010", -- 12
		       "00000000000010000000000000000000" when "10011", -- 13
		       "00000000000100000000000000000000" when "10100", -- 14
		       "00000000001000000000000000000000" when "10101", -- 15
		       "00000000010000000000000000000000" when "10110", -- 16
		       "00000000100000000000000000000000" when "10111", -- 17
		       "00000001000000000000000000000000" when "11000", -- 18
		       "00000010000000000000000000000000" when "11001", -- 19
		       "00000100000000000000000000000000" when "11010", -- 1A
		       "00001000000000000000000000000000" when "11011", -- 1B
		       "00010000000000000000000000000000" when "11100", -- 1C
		       "00100000000000000000000000000000" when "11101", -- 1D
		       "01000000000000000000000000000000" when "11110", -- 1E
		       "10000000000000000000000000000000" when "11111", -- 1F
		       "00000000000000000000000000000000" when others;  -- other
end dataflow;
