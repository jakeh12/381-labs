jhladik@Jakubs-MacBook-Pro.local.2533